module divide64x16x51x16 (reset, A, B, Qout, clk);

	input reset;
    input[64 - 1:0] A; 
    input[51 - 1:0] B; 
    output[16 - 1:0] Qout; 
    reg[16 - 1:0] Qout;
    input clk; 

    reg[64 + 16 - 1:0] c0; 
    reg[64 + 16 - 1:0] c1; 
    reg[64 + 16 - 1:0] c2; 
    reg[64 + 16 - 1:0] c3; 
    reg[64 + 16 - 1:0] c4; 
    reg[64 + 16 - 1:0] c5; 
    reg[64 + 16 - 1:0] c6; 
    reg[64 + 16 - 1:0] c7; 
    reg[64 + 16 - 1:0] c8; 
    reg[64 + 16 - 1:0] c9; 
    reg[64 + 16 - 1:0] c10; 
    reg[64 + 16 - 1:0] c11; 
    reg[64 + 16 - 1:0] c12; 
    reg[64 + 16 - 1:0] c13; 
    reg[64 + 16 - 1:0] c14; 
    reg[64 + 16 - 1:0] c15; 

    reg[16 - 1:0] q0; 
	reg[16 - 1:0] q1; 
    reg[16 - 1:0] q2; 
    reg[16 - 1:0] q3; 
    reg[16 - 1:0] q4; 
    reg[16 - 1:0] q5; 
    reg[16 - 1:0] q6; 
    reg[16 - 1:0] q7; 
    reg[16 - 1:0] q8; 
    reg[16 - 1:0] q9; 
    reg[16 - 1:0] q10; 
	reg[16 - 1:0] q11; 
    reg[16 - 1:0] q12; 
    reg[16 - 1:0] q13; 
    reg[16 - 1:0] q14; 
    reg[16 - 1:0] q15; 

    reg[51 - 1:0] bp0; 
    reg[51 - 1:0] bp1; 
    reg[51 - 1:0] bp2; 
    reg[51 - 1:0] bp3; 
    reg[51 - 1:0] bp4; 
    reg[51 - 1:0] bp5; 
    reg[51 - 1:0] bp6; 
    reg[51 - 1:0] bp7; 
    reg[51 - 1:0] bp8; 
    reg[51 - 1:0] bp9; 
    reg[51 - 1:0] bp10; 
    reg[51 - 1:0] bp11; 
    reg[51 - 1:0] bp12; 
    reg[51 - 1:0] bp13; 
    reg[51 - 1:0] bp14; 
    reg[51 - 1:0] bp15; 

    always @(posedge clk or negedge reset)
    begin
	if (reset == 1'b0)
	begin

    c0 <= 0; 
    c1 <= 0; 
    c2 <= 0; 
    c3 <= 0; 
    c4 <= 0; 
    c5 <= 0; 
    c6 <= 0; 
    c7 <= 0; 
    c8 <= 0; 
    c9 <= 0; 
    c10 <= 0; 
    c11 <= 0; 
    c12 <= 0; 
    c13 <= 0; 
    c14 <= 0; 
    c15 <= 0; 
        q0 <= 0; 
	q1 <= 0; 
    q2 <= 0; 
    q3 <= 0; 
    q4 <= 0; 
    q5 <= 0; 
    q6 <= 0; 
    q7 <= 0; 
    q8 <= 0; 
    q9 <= 0; 
    q10 <= 0; 
	q11 <= 0; 
    q12 <= 0; 
    q13 <= 0; 
    q14 <= 0; 
        bp0 <= 0; 
    bp1 <= 0; 
    bp2 <= 0; 
    bp3 <= 0; 
    bp4 <= 0; 
    bp5 <= 0; 
    bp6 <= 0; 
    bp7 <= 0; 
    bp8 <= 0; 
    bp9 <= 0; 
    bp10 <= 0; 
    bp11 <= 0; 
    bp12 <= 0; 
    bp13 <= 0; 
    bp14 <= 0; 
    bp15 <= 0; 
   	end
	else
	begin


    c0[64 + 16 - 1:16] <= A ;
    c0[16 - 1:0] <= 0;
    q0 <= 0;
    bp0 <= B ;
	bp1 <= bp0 ;
    bp2 <= bp1 ;
    bp3 <= bp2 ;
    bp4 <= bp3 ;
    bp5 <= bp4 ;
    bp6 <= bp5 ;
    bp7 <= bp6 ;
    bp8 <= bp7 ;
    bp9 <= bp8 ;
    bp10 <= bp9 ;
    bp11 <= bp10 ;
    bp12 <= bp11 ;
    bp13 <= bp12 ;
    bp14 <= bp13 ;
    bp15 <= bp14 ;


		if (c0[64 + 16 - 1:16 - 1 - 0] >= bp0[47:0] )
		begin
			q1 <= {q0[16-2:0] , 1'b1}; 
 			c1 <= {(c0[64+16-1:16-1-0] - bp0[47:0]), c0[16-0-2:0]} ; 
		end
		else
		begin
			q1 <= {q0[16-2:0], 1'b0} ; 
			c1 <= c0 ; 
		end
		if (c1[64 + 16 - 1:16 - 1 - 1] >= bp1[47:0] )
		begin
			q2 <= {q1[16-2:0] , 1'b1}; 
 			c2 <= {(c1[64+16-1:16-1-1] - bp1[47:0]), c1[16-1-2:0]} ; 
		end
		else
		begin
			q2 <= {q1[16-2:0], 1'b0} ; 
			c2 <= c1 ; 
		end
		if (c2[64 + 16 - 1:16 - 1 - 2] >= bp2[47:0] )
		begin
			q3 <= {q2[16-2:0] , 1'b1}; 
 			c3 <= {(c2[64+16-1:16-1-2] - bp2[47:0]), c2[16-2-2:0]} ; 
		end
		else
		begin
			q3 <= {q2[16-2:0], 1'b0} ; 
			c3 <= c2 ; 
		end
		if (c3[64 + 16 - 1:16 - 1 - 3] >= bp3[47:0] )
		begin
			q4 <= {q3[16-2:0] , 1'b1}; 
 			c4 <= {(c3[64+16-1:16-1-3] - bp3[47:0]), c3[16-3-2:0]} ; 
		end
		else
		begin
			q4 <= {q3[16-2:0], 1'b0} ; 
			c4 <= c3 ; 
		end
		if (c4[64 + 16 - 1:16 - 1 - 4] >= bp4[47:0] )
		begin
			q5 <= {q4[16-2:0] , 1'b1}; 
 			c5 <= {(c4[64+16-1:16-1-4] - bp4[47:0]), c4[16-4-2:0]} ; 
		end
		else
		begin
			q5 <= {q4[16-2:0], 1'b0} ; 
			c5 <= c4 ; 
		end
		if (c5[64 + 16 - 1:16 - 1 - 5] >= bp5[47:0] )
		begin
			q6 <= {q5[16-2:0] , 1'b1}; 
 			c6 <= {(c5[64+16-1:16-1-5] - bp5[47:0]), c5[16-5-2:0]} ; 
		end
		else
		begin
			q6 <= {q5[16-2:0], 1'b0} ; 
			c6 <= c5 ; 
		end
		if (c6[64 + 16 - 1:16 - 1 - 6] >= bp6[47:0] )
		begin
			q7 <= {q6[16-2:0] , 1'b1}; 
 			c7 <= {(c6[64+16-1:16-1-6] - bp6[47:0]), c6[16-6-2:0]} ; 
		end
		else
		begin
			q7 <= {q6[16-2:0], 1'b0} ; 
			c7 <= c6 ; 
		end
		if (c7[64 + 16 - 1:16 - 1 - 7] >= bp7[47:0] )
		begin
			q8 <= {q7[16-2:0] , 1'b1}; 
 			c8 <= {(c7[64+16-1:16-1-7] - bp7[47:0]), c7[16-7-2:0]} ; 
		end
		else
		begin
			q8 <= {q7[16-2:0], 1'b0} ; 
			c8 <= c7 ; 
		end
		if (c8[64 + 16 - 1:16 - 1 - 8] >= bp8[47:0] )
		begin
			q9 <= {q8[16-2:0] , 1'b1}; 
 			c9 <= {(c8[64+16-1:16-1-8] - bp8[47:0]), c8[16-8-2:0]} ; 
		end
		else
		begin
			q9 <= {q8[16-2:0], 1'b0} ; 
			c9 <= c8 ; 
		end
		if (c9[64 + 16 - 1:16 - 1 - 9] >= bp9[47:0] )
		begin
			q10 <= {q9[16-2:0] , 1'b1}; 
 			c10 <= {(c9[64+16-1:16-1-9] - bp9[47:0]), c9[16-9-2:0]} ; 
		end
		else
		begin
			q10 <= {q9[16-2:0], 1'b0} ; 
			c10 <= c9 ; 
		end
		if (c10[64 + 16 - 1:16 - 1 - 10] >= bp10[47:0] )
		begin
			q11 <= {q10[16-2:0] , 1'b1}; 
 			c11 <= {(c10[64+16-1:16-1-10] - bp10[47:0]), c10[16-10-2:0]} ; 
		end
		else
		begin
			q11 <= {q10[16-2:0], 1'b0} ; 
			c11 <= c10 ; 
		end

		if (c11[64 + 16 - 1:16 - 1 - 11] >= bp11[47:0] )
		begin
			q12 <= {q11[16-2:0] , 1'b1}; 
 			c12 <= {(c11[64+16-1:16-1-11] - bp11[47:0]), c11[16-11-2:0]} ; 
		end
		else
		begin
			q12 <= {q11[16-2:0], 1'b0} ; 
			c12 <= c11 ; 
		end
		if (c12[64 + 16 - 1:16 - 1 - 12] >= bp12[47:0] )
		begin
			q13 <= {q12[16-2:0] , 1'b1}; 
 			c13 <= {(c12[64+16-1:16-1-12] - bp12[47:0]), c12[16-12-2:0]} ; 
		end
		else
		begin
			q13 <= {q12[16-2:0], 1'b0} ; 
			c13 <= c12 ; 
		end
		if (c13[64 + 16 - 1:16 - 1 - 13] >= bp13[47:0] )
		begin
			q14 <= {q13[16-2:0] , 1'b1}; 
 			c14 <= {(c13[64+16-1:16-1-13] - bp13[47:0]), c13[16-13-2:0]} ; 
		end
		else
		begin
			q14 <= {q13[16-2:0], 1'b0} ; 
			c14 <= c13 ; 
		end
		if (c14[64 + 16 - 1:16 - 1 - 14] >= bp14[47:0] )
		begin
			q15 <= {q14[16-2:0] , 1'b1}; 
 			c15 <= {(c14[64+16-1:16-1-14] - bp14[47:0]), c14[16-14-2:0]} ; 
		end
		else
		begin
			q15 <= {q14[16-2:0], 1'b0} ; 
			c15 <= c14 ; 
		end

          if (c15 >= bp15 )
          begin
             Qout <= {q15[16-2:0], 1'b1} ; 
          end
          else
          begin
             Qout <= {q15[16-2:0], 1'b0} ; 
          end 
	end
    end 
 endmodule