module divide64x32x51x18 (reset, A, B, Qout, clk);

	input reset;
    input[64 - 1:0] A; 
    input[51 - 1:0] B; 
    output[32 - 1:0] Qout; 
    reg[32 - 1:0] Qout;
    input clk; 

    reg[64 + 15 - 1:0] c0; 
    reg[64 + 15 - 1:0] c1; 
    reg[64 + 15 - 1:0] c2; 
    reg[64 + 15 - 1:0] c3; 
    reg[64 + 15 - 1:0] c4; 
    reg[64 + 15 - 1:0] c5; 
    reg[64 + 15 - 1:0] c6; 
    reg[64 + 15 - 1:0] c7; 
    reg[64 + 15 - 1:0] c8; 
    reg[64 + 15 - 1:0] c9; 
    reg[64 + 15 - 1:0] c10; 
    reg[64 + 15 - 1:0] c11; 
    reg[64 + 15 - 1:0] c12; 
    reg[64 + 15 - 1:0] c13; 
    reg[64 + 15 - 1:0] c14; 
    reg[64 + 15 - 1:0] c15; 
    reg[64 + 15 - 1:0] c16; 
    reg[64 + 15 - 1:0] c17; 
    reg[64 + 15 - 1:0] c18; 
    reg[64 + 15 - 1:0] c19; 
    reg[64 + 15 - 1:0] c20; 
    reg[64 + 15 - 1:0] c21; 
    reg[64 + 15 - 1:0] c22; 
    reg[64 + 15 - 1:0] c23; 
    reg[64 + 15 - 1:0] c24; 
    reg[64 + 15 - 1:0] c25; 
    reg[64 + 15 - 1:0] c26; 
    reg[64 + 15 - 1:0] c27; 
    reg[64 + 15 - 1:0] c28; 
    reg[64 + 15 - 1:0] c29; 
    reg[64 + 15 - 1:0] c30; 
    reg[64 + 15 - 1:0] c31; 

    reg[32 - 1:0] q0; 
	reg[32 - 1:0] q1; 
    reg[32 - 1:0] q2; 
    reg[32 - 1:0] q3; 
    reg[32 - 1:0] q4; 
    reg[32 - 1:0] q5; 
    reg[32 - 1:0] q6; 
    reg[32 - 1:0] q7; 
    reg[32 - 1:0] q8; 
    reg[32 - 1:0] q9; 
    reg[32 - 1:0] q10; 
	reg[32 - 1:0] q11; 
    reg[32 - 1:0] q12; 
    reg[32 - 1:0] q13; 
    reg[32 - 1:0] q14; 
    reg[32 - 1:0] q15; 
    reg[32 - 1:0] q16; 
    reg[32 - 1:0] q17; 
    reg[32 - 1:0] q18; 
    reg[32 - 1:0] q19; 
    reg[32 - 1:0] q20; 
	reg[32 - 1:0] q21; 
    reg[32 - 1:0] q22; 
    reg[32 - 1:0] q23; 
    reg[32 - 1:0] q24; 
    reg[32 - 1:0] q25; 
    reg[32 - 1:0] q26; 
    reg[32 - 1:0] q27; 
    reg[32 - 1:0] q28; 
    reg[32 - 1:0] q29; 
    reg[32 - 1:0] q30; 
    reg[32 - 1:0] q31; 

    reg[51 - 1:0] bp0; 
    reg[51 - 1:0] bp1; 
    reg[51 - 1:0] bp2; 
    reg[51 - 1:0] bp3; 
    reg[51 - 1:0] bp4; 
    reg[51 - 1:0] bp5; 
    reg[51 - 1:0] bp6; 
    reg[51 - 1:0] bp7; 
    reg[51 - 1:0] bp8; 
    reg[51 - 1:0] bp9; 
    reg[51 - 1:0] bp10; 
    reg[51 - 1:0] bp11; 
    reg[51 - 1:0] bp12; 
    reg[51 - 1:0] bp13; 
    reg[51 - 1:0] bp14; 
    reg[51 - 1:0] bp15; 
    reg[51 - 1:0] bp16; 
    reg[51 - 1:0] bp17; 
    reg[51 - 1:0] bp18; 
    reg[51 - 1:0] bp19; 
    reg[51 - 1:0] bp20; 
    reg[51 - 1:0] bp21; 
    reg[51 - 1:0] bp22; 
    reg[51 - 1:0] bp23; 
    reg[51 - 1:0] bp24; 
    reg[51 - 1:0] bp25; 
    reg[51 - 1:0] bp26; 
    reg[51 - 1:0] bp27; 
    reg[51 - 1:0] bp28; 
    reg[51 - 1:0] bp29; 
    reg[51 - 1:0] bp30; 
    reg[51 - 1:0] bp31; 

    reg [64 + 15 - 1:0] c_xhdl;

	always @(posedge clk or negedge reset)
    begin
	if (reset == 1'b0)
	begin

    c0 <= 0; 
    c1 <= 0; 
    c2 <= 0; 
    c3 <= 0; 
    c4 <= 0; 
    c5 <= 0; 
    c6 <= 0; 
    c7 <= 0; 
    c8 <= 0; 
    c9 <= 0; 
    c10 <= 0; 
    c11 <= 0; 
    c12 <= 0; 
    c13 <= 0; 
    c14 <= 0; 
    c15 <= 0; 
    c16 <= 0; 
    c17 <= 0; 
    c18 <= 0; 
    c19 <= 0; 
    c20 <= 0; 
    c21 <= 0; 
    c22 <= 0; 
    c23 <= 0; 
    c24 <= 0; 
    c25 <= 0; 
    c26 <= 0; 
    c27 <= 0; 
    c28 <= 0; 
    c29 <= 0; 
    c30 <= 0; 
    c31 <= 0; 

    q0 <= 0; 
	q1 <= 0; 
    q2 <= 0; 
    q3 <= 0; 
    q4 <= 0; 
    q5 <= 0; 
    q6 <= 0; 
    q7 <= 0; 
    q8 <= 0; 
    q9 <= 0; 
    q10 <= 0; 
	q11 <= 0; 
    q12 <= 0; 
    q13 <= 0; 
    q14 <= 0; 
    q15 <= 0; 
    q16 <= 0; 
    q17 <= 0; 
    q18 <= 0; 
    q19 <= 0; 
    q20 <= 0; 
	q21 <= 0; 
    q22 <= 0; 
    q23 <= 0; 
    q24 <= 0; 
    q25 <= 0; 
    q26 <= 0; 
    q27 <= 0; 
    q28 <= 0; 
    q29 <= 0; 
    q30 <= 0; 
    q31 <= 0; 

    bp0 <= 0; 
    bp1 <= 0; 
    bp2 <= 0; 
    bp3 <= 0; 
    bp4 <= 0; 
    bp5 <= 0; 
    bp6 <= 0; 
    bp7 <= 0; 
    bp8 <= 0; 
    bp9 <= 0; 
    bp10 <= 0; 
    bp11 <= 0; 
    bp12 <= 0; 
    bp13 <= 0; 
    bp14 <= 0; 
    bp15 <= 0; 
    bp16 <= 0; 
    bp17 <= 0; 
    bp18 <= 0; 
    bp19 <= 0; 
    bp20 <= 0; 
    bp21 <= 0; 
    bp22 <= 0; 
    bp23 <= 0; 
    bp24 <= 0; 
    bp25 <= 0; 
    bp26 <= 0; 
    bp27 <= 0; 
    bp28 <= 0; 
    bp29 <= 0; 
    bp30 <= 0; 
    bp31 <= 0; 

	end
	else
	begin

    c0[64 + 15 - 1:15] <= A ;
    c0[15 - 1:0] <= 0;
    q0 <= 0;
    bp0 <= B ;
    bp1 <= bp0 ;
    bp2 <= bp1 ;
    bp3 <= bp2 ;
    bp4 <= bp3 ;
    bp5 <= bp4 ;
    bp6 <= bp5 ;
    bp7 <= bp6 ;
    bp8 <= bp7 ;
    bp9 <= bp8 ;
    bp10 <= bp9 ;
    bp11 <= bp10 ;
    bp12 <= bp11 ;
    bp13 <= bp12 ;
    bp14 <= bp13 ;
    bp15 <= bp14 ;
    bp16 <= bp15 ;
    bp17 <= bp16 ;
    bp18 <= bp17 ;
    bp19 <= bp18 ;
    bp20 <= bp19 ;
    bp21 <= bp20 ;
    bp22 <= bp21 ;
    bp23 <= bp22 ;
    bp24 <= bp23 ;
    bp25 <= bp24 ;
    bp26 <= bp25 ;
    bp27 <= bp26 ;
    bp28 <= bp27 ;
    bp29 <= bp28 ;
    bp30 <= bp29 ;
    bp31 <= bp30 ;

		if (c0[64 + 15 - 1:32 - 1 - 0] >= bp0[47:0] )
		begin
			q1 <= {q0[32-2:0] , 1'b1}; 
 			c1 <= {(c0[64+15-1:32-1-0] - bp0[47:0]), c0[32-0-2:0]} ; 
		end
		else
		begin
			q1 <= {q0[32-2:0], 1'b0} ; 
			c1 <= c0 ; 
		end
		if (c1[64 + 15 - 1:32 - 1 - 1] >= bp1[47:0] )
		begin
			q2 <= {q1[32-2:0] , 1'b1}; 
 			c2 <= {(c1[64+15-1:32-1-1] - bp1[47:0]), c1[32-1-2:0]} ; 
		end
		else
		begin
			q2 <= {q1[32-2:0], 1'b0} ; 
			c2 <= c1 ; 
		end
		if (c2[64 + 15 - 1:32 - 1 - 2] >= bp2[47:0] )
		begin
			q3 <= {q2[32-2:0] , 1'b1}; 
 			c3 <= {(c2[64+15-1:32-1-2] - bp2[47:0]), c2[32-2-2:0]} ; 
		end
		else
		begin
			q3 <= {q2[32-2:0], 1'b0} ; 
			c3 <= c2 ; 
		end
		if (c3[64 + 15 - 1:32 - 1 - 3] >= bp3[47:0] )
		begin
			q4 <= {q3[32-2:0] , 1'b1}; 
 			c4 <= {(c3[64+15-1:32-1-3] - bp3[47:0]), c3[32-3-2:0]} ; 
		end
		else
		begin
			q4 <= {q3[32-2:0], 1'b0} ; 
			c4 <= c3 ; 
		end
		if (c4[64 + 15 - 1:32 - 1 - 4] >= bp4[47:0] )
		begin
			q5 <= {q4[32-2:0] , 1'b1}; 
 			c5 <= {(c4[64+15-1:32-1-4] - bp4[47:0]), c4[32-4-2:0]} ; 
		end
		else
		begin
			q5 <= {q4[32-2:0], 1'b0} ; 
			c5 <= c4 ; 
		end
		if (c5[64 + 15 - 1:32 - 1 - 5] >= bp5[47:0] )
		begin
			q6 <= {q5[32-2:0] , 1'b1}; 
 			c6 <= {(c5[64+15-1:32-1-5] - bp5[47:0]), c5[32-5-2:0]} ; 
		end
		else
		begin
			q6 <= {q5[32-2:0], 1'b0} ; 
			c6 <= c5 ; 
		end
		if (c6[64 + 15 - 1:32 - 1 - 6] >= bp6[47:0] )
		begin
			q7 <= {q6[32-2:0] , 1'b1}; 
 			c7 <= {(c6[64+15-1:32-1-6] - bp6[47:0]), c6[32-6-2:0]} ; 
		end
		else
		begin
			q7 <= {q6[32-2:0], 1'b0} ; 
			c7 <= c6 ; 
		end
		if (c7[64 + 15 - 1:32 - 1 - 7] >= bp7[47:0] )
		begin
			q8 <= {q7[32-2:0] , 1'b1}; 
 			c8 <= {(c7[64+15-1:32-1-7] - bp7[47:0]), c7[32-7-2:0]} ; 
		end
		else
		begin
			q8 <= {q7[32-2:0], 1'b0} ; 
			c8 <= c7 ; 
		end
		if (c8[64 + 15 - 1:32 - 1 - 8] >= bp8[47:0] )
		begin
			q9 <= {q8[32-2:0] , 1'b1}; 
 			c9 <= {(c8[64+15-1:32-1-8] - bp8[47:0]), c8[32-8-2:0]} ; 
		end
		else
		begin
			q9 <= {q8[32-2:0], 1'b0} ; 
			c9 <= c8 ; 
		end
		if (c9[64 + 15 - 1:32 - 1 - 9] >= bp9[47:0] )
		begin
			q10 <= {q9[32-2:0] , 1'b1}; 
 			c10 <= {(c9[64+15-1:32-1-9] - bp9[47:0]), c9[32-9-2:0]} ; 
		end
		else
		begin
			q10 <= {q9[32-2:0], 1'b0} ; 
			c10 <= c9 ; 
		end
		if (c10[64 + 15 - 1:32 - 1 - 10] >= bp10[47:0] )
		begin
			q11 <= {q10[32-2:0] , 1'b1}; 
 			c11 <= {(c10[64+15-1:32-1-10] - bp10[47:0]), c10[32-10-2:0]} ; 
		end
		else
		begin
			q11 <= {q10[32-2:0], 1'b0} ; 
			c11 <= c10 ; 
		end

		if (c11[64 + 15 - 1:32 - 1 - 11] >= bp11[47:0] )
		begin
			q12 <= {q11[32-2:0] , 1'b1}; 
 			c12 <= {(c11[64+15-1:32-1-11] - bp11[47:0]), c11[32-11-2:0]} ; 
		end
		else
		begin
			q12 <= {q11[32-2:0], 1'b0} ; 
			c12 <= c11 ; 
		end
		if (c12[64 + 15 - 1:32 - 1 - 12] >= bp12[47:0] )
		begin
			q13 <= {q12[32-2:0] , 1'b1}; 
 			c13 <= {(c12[64+15-1:32-1-12] - bp12[47:0]), c12[32-12-2:0]} ; 
		end
		else
		begin
			q13 <= {q12[32-2:0], 1'b0} ; 
			c13 <= c12 ; 
		end
		if (c13[64 + 15 - 1:32 - 1 - 13] >= bp13[47:0] )
		begin
			q14 <= {q13[32-2:0] , 1'b1}; 
 			c14 <= {(c13[64+15-1:32-1-13] - bp13[47:0]), c13[32-13-2:0]} ; 
		end
		else
		begin
			q14 <= {q13[32-2:0], 1'b0} ; 
			c14 <= c13 ; 
		end
		if (c14[64 + 15 - 1:32 - 1 - 14] >= bp14[47:0] )
		begin
			q15 <= {q14[32-2:0] , 1'b1}; 
 			c15 <= {(c14[64+15-1:32-1-14] - bp14[47:0]), c14[32-14-2:0]} ; 
		end
		else
		begin
			q15 <= {q14[32-2:0], 1'b0} ; 
			c15 <= c14 ; 
		end
		if (c15[64 + 15 - 1:32 - 1 - 15] >= bp15[47:0] )
		begin
			q16 <= {q15[32-2:0] , 1'b1}; 
 			c16 <= {(c15[64+15-1:32-1-15] - bp15[47:0]), c15[32-15-2:0]} ; 
		end
		else
		begin
			q16 <= {q15[32-2:0], 1'b0} ; 
			c16 <= c15 ; 
		end
		if (c16[64 + 15 - 1:32 - 1 - 16] >= bp16[47:0] )
		begin
			q17 <= {q16[32-2:0] , 1'b1}; 
 			c17 <= {(c16[64+15-1:32-1-16] - bp16[47:0]), c16[32-16-2:0]} ; 
		end
		else
		begin
			q17 <= {q16[32-2:0], 1'b0} ; 
			c17 <= c16 ; 
		end
		if (c17[64 + 15 - 1:32 - 1 - 17] >= bp17[47:0] )
		begin
			q18 <= {q17[32-2:0] , 1'b1}; 
 			c18 <= {(c17[64+15-1:32-1-17] - bp17[47:0]), c17[32-17-2:0]} ; 
		end
		else
		begin
			q18 <= {q17[32-2:0], 1'b0} ; 
			c18 <= c17 ; 
		end
		if (c18[64 + 15 - 1:32 - 1 - 18] >= bp18[47:0] )
		begin
			q19 <= {q18[32-2:0] , 1'b1}; 
 			c19 <= {(c18[64+15-1:32-1-18] - bp18[47:0]), c18[32-18-2:0]} ; 
		end
		else
		begin
			q19 <= {q18[32-2:0], 1'b0} ; 
			c19 <= c18 ; 
		end
		if (c19[64 + 15 - 1:32 - 1 - 19] >= bp19[47:0] )
		begin
			q20 <= {q19[32-2:0] , 1'b1}; 
 			c20 <= {(c19[64+15-1:32-1-19] - bp19[47:0]), c19[32-19-2:0]} ; 
		end
		else
		begin
			q20 <= {q19[32-2:0], 1'b0} ; 
			c20 <= c19 ; 
		end

		if (c20[64 + 15 - 1:32 - 1 - 20] >= bp20[47:0] )
		begin
			q21 <= {q20[32-2:0] , 1'b1}; 
 			c21 <= {(c20[64+15-1:32-1-20] - bp20[47:0]), c20[32-20-2:0]} ; 
		end
		else
		begin
			q21 <= {q20[32-2:0], 1'b0} ; 
			c21 <= c20 ; 
		end
		if (c21[64 + 15 - 1:32 - 1 - 21] >= bp21[47:0] )
		begin
			q22 <= {q21[32-2:0] , 1'b1}; 
 			c22 <= {(c21[64+15-1:32-1-21] - bp21[47:0]), c21[32-21-2:0]} ; 
		end
		else
		begin
			q22 <= {q21[32-2:0], 1'b0} ; 
			c22 <= c21 ; 
		end
		if (c22[64 + 15 - 1:32 - 1 - 22] >= bp22[47:0] )
		begin
			q23 <= {q22[32-2:0] , 1'b1}; 
 			c23 <= {(c22[64+15-1:32-1-22] - bp22[47:0]), c22[32-22-2:0]} ; 
		end
		else
		begin
			q23 <= {q22[32-2:0], 1'b0} ; 
			c23 <= c22; 
		end
		if (c23[64 + 15 - 1:32 - 1 - 23] >= bp23[47:0] )
		begin
			q24 <= {q23[32-2:0] , 1'b1}; 
 			c24 <= {(c23[64+15-1:32-1-23] - bp23[47:0]), c23[32-23-2:0]} ; 
		end
		else
		begin
			q24 <= {q23[32-2:0], 1'b0} ; 
			c24 <= c23 ; 
		end
		if (c24[64 + 15 - 1:32 - 1 - 24] >= bp24[47:0] )
		begin
			q25 <= {q24[32-2:0] , 1'b1}; 
 			c25 <= {(c24[64+15-1:32-1-24] - bp24[47:0]), c24[32-24-2:0]} ; 
		end
		else
		begin
			q25 <= {q24[32-2:0], 1'b0} ; 
			c25 <= c24 ; 
		end
		if (c25[64 + 15 - 1:32 - 1 - 25] >= bp25[47:0] )
		begin
			q26 <= {q25[32-2:0] , 1'b1}; 
 			c26 <= {(c25[64+15-1:32-1-25] - bp25[47:0]), c25[32-25-2:0]} ; 
		end
		else
		begin
			q26 <= {q25[32-2:0], 1'b0} ; 
			c26 <= c25 ; 
		end
		if (c26[64 + 15 - 1:32 - 1 - 26] >= bp26[47:0] )
		begin
			q27 <= {q26[32-2:0] , 1'b1}; 
 			c27 <= {(c26[64+15-1:32-1-26] - bp26[47:0]), c26[32-26-2:0]} ; 
		end
		else
		begin
			q27 <= {q26[32-2:0], 1'b0} ; 
			c27 <= c26 ; 
		end
		if (c27[64 + 15 - 1:32 - 1 - 27] >= bp27[47:0] )
		begin
			q28 <= {q27[32-2:0] , 1'b1}; 
 			c28 <= {(c27[64+15-1:32-1-27] - bp27[47:0]), c27[32-27-2:0]} ; 
		end
		else
		begin
			q28 <= {q27[32-2:0], 1'b0} ; 
			c28 <= c27 ; 
		end
		if (c28[64 + 15 - 1:32 - 1 - 29] >= bp28[47:0] )
		begin
			q29 <= {q28[32-2:0] , 1'b1}; 
 			c29 <= {(c28[64+15-1:32-1-29] - bp28[47:0]), c28[32-29-2:0]} ; 
		end
		else
		begin
			q29 <= {q28[32-2:0], 1'b0} ; 
			c29 <= c28 ; 
		end
		if (c29[64 + 15 - 1:32 - 1 - 29] >= bp29[47:0] )
		begin
			q30 <= {q29[32-2:0] , 1'b1}; 
 			c30 <= {(c29[64+15-1:32-1-29] - bp29[47:0]), c29[32-29-2:0]} ; 
		end
		else
		begin
			q30 <= {q29[32-2:0], 1'b0} ; 
			c30 <= c29 ; 
		end
		if (c30[64 + 15 - 1:32 - 1 - 30] >= bp30[47:0] )
		begin
			q31 <= {q30[32-2:0] , 1'b1}; 
 			c31 <= {(c30[64+15-1:32-1-30] - bp30[47:0]), c30[32-30-2:0]} ; 
		end
		else
		begin
			q31 <= {q30[32-2:0], 1'b0} ; 
			c31 <= c30 ; 
		end

          if (c31 >= bp31 )
          begin
             Qout <= {q31[32-2:0], 1'b1} ; 
          end
          else
          begin
             Qout <= {q31[32-2:0], 1'b0} ; 
          end 
	end
    end 
 endmodule