module Sorter (clk, rst_n, guard, value, reg_0);
integer index; // Used for initialisations
input clk;
input rst_n;
output guard;
output [63:0] value;
// state declarations
input [63:0] reg_0;
// bindings 
wire  wire0 = 0'b0;
wire  wire1 = 1'b1;
wire  wire2 = 1'b0;
wire [63:0] wire3 = reg_0;
wire [31:0] wire4 = wire3[31:0];
wire [31:0] wire5 = wire3[63:32];
wire [31:0] wire6 = wire5[31:0];
wire [15:0] wire7 = wire4[15:0];
wire [15:0] wire8 = wire4[31:16];
wire [15:0] wire9 = wire8[15:0];
wire [7:0] wire10 = wire7[7:0];
wire [7:0] wire11 = wire7[15:8];
wire [7:0] wire12 = wire11[7:0];
wire [3:0] wire13 = wire10[3:0];
wire [3:0] wire14 = wire10[7:4];
wire [3:0] wire15 = wire14[3:0];
wire [3:0] wire16 = wire12[3:0];
wire [3:0] wire17 = wire12[7:4];
wire [3:0] wire18 = wire17[3:0];
wire [7:0] wire19 = wire9[7:0];
wire [7:0] wire20 = wire9[15:8];
wire [7:0] wire21 = wire20[7:0];
wire [3:0] wire22 = wire19[3:0];
wire [3:0] wire23 = wire19[7:4];
wire [3:0] wire24 = wire23[3:0];
wire [3:0] wire25 = wire21[3:0];
wire [3:0] wire26 = wire21[7:4];
wire [3:0] wire27 = wire26[3:0];
wire [15:0] wire28 = wire6[15:0];
wire [15:0] wire29 = wire6[31:16];
wire [15:0] wire30 = wire29[15:0];
wire [7:0] wire31 = wire28[7:0];
wire [7:0] wire32 = wire28[15:8];
wire [7:0] wire33 = wire32[7:0];
wire [3:0] wire34 = wire31[3:0];
wire [3:0] wire35 = wire31[7:4];
wire [3:0] wire36 = wire35[3:0];
wire [3:0] wire37 = wire33[3:0];
wire [3:0] wire38 = wire33[7:4];
wire [3:0] wire39 = wire38[3:0];
wire [7:0] wire40 = wire30[7:0];
wire [7:0] wire41 = wire30[15:8];
wire [7:0] wire42 = wire41[7:0];
wire [3:0] wire43 = wire40[3:0];
wire [3:0] wire44 = wire40[7:4];
wire [3:0] wire45 = wire44[3:0];
wire [3:0] wire46 = wire42[3:0];
wire [3:0] wire47 = wire42[7:4];
wire [3:0] wire48 = wire47[3:0];
wire [7:0] wire49 = {wire13, wire15};
wire [3:0] wire50 = wire49[7:4];
wire  wire51 = wire13 <= wire15;
wire [3:0] wire52 = wire51 ? wire13 : wire15;
wire [3:0] wire53 = wire51 ? wire15 : wire13;
wire [7:0] wire54 = {wire52, wire53};
wire [3:0] wire55 = wire54[7:4];
wire [7:0] wire56 = {wire16, wire18};
wire [3:0] wire57 = wire56[7:4];
wire  wire58 = wire16 <= wire18;
wire [3:0] wire59 = wire58 ? wire16 : wire18;
wire [3:0] wire60 = wire58 ? wire18 : wire16;
wire [7:0] wire61 = {wire59, wire60};
wire [3:0] wire62 = wire61[7:4];
wire [7:0] wire63 = {wire60, wire59};
wire [15:0] wire64 = {wire54, wire63};
wire [7:0] wire65 = wire64[15:8];
wire [3:0] wire66 = wire63[7:4];
wire  wire67 = wire52 <= wire60;
wire [3:0] wire68 = wire67 ? wire52 : wire60;
wire [3:0] wire69 = wire67 ? wire60 : wire52;
wire [7:0] wire70 = {wire68, wire69};
wire [3:0] wire71 = wire70[7:4];
wire  wire72 = wire53 <= wire59;
wire [3:0] wire73 = wire72 ? wire53 : wire59;
wire [3:0] wire74 = wire72 ? wire59 : wire53;
wire [7:0] wire75 = {wire73, wire74};
wire [3:0] wire76 = wire75[7:4];
wire [7:0] wire77 = {wire68, wire73};
wire [7:0] wire78 = {wire69, wire74};
wire [15:0] wire79 = {wire77, wire78};
wire [7:0] wire80 = wire79[15:8];
wire [3:0] wire81 = wire77[7:4];
wire  wire82 = wire68 <= wire73;
wire [3:0] wire83 = wire82 ? wire68 : wire73;
wire [3:0] wire84 = wire82 ? wire73 : wire68;
wire [7:0] wire85 = {wire83, wire84};
wire [3:0] wire86 = wire85[7:4];
wire  wire87 = wire69 <= wire74;
wire [3:0] wire88 = wire87 ? wire69 : wire74;
wire [3:0] wire89 = wire87 ? wire74 : wire69;
wire [7:0] wire90 = {wire88, wire89};
wire [3:0] wire91 = wire90[7:4];
wire [15:0] wire92 = {wire85, wire90};
wire [7:0] wire93 = {wire22, wire24};
wire [3:0] wire94 = wire93[7:4];
wire  wire95 = wire22 <= wire24;
wire [3:0] wire96 = wire95 ? wire22 : wire24;
wire [3:0] wire97 = wire95 ? wire24 : wire22;
wire [7:0] wire98 = {wire96, wire97};
wire [3:0] wire99 = wire98[7:4];
wire [7:0] wire100 = {wire25, wire27};
wire [3:0] wire101 = wire100[7:4];
wire  wire102 = wire25 <= wire27;
wire [3:0] wire103 = wire102 ? wire25 : wire27;
wire [3:0] wire104 = wire102 ? wire27 : wire25;
wire [7:0] wire105 = {wire103, wire104};
wire [3:0] wire106 = wire105[7:4];
wire [7:0] wire107 = {wire104, wire103};
wire [15:0] wire108 = {wire98, wire107};
wire [7:0] wire109 = wire108[15:8];
wire [3:0] wire110 = wire107[7:4];
wire  wire111 = wire96 <= wire104;
wire [3:0] wire112 = wire111 ? wire96 : wire104;
wire [3:0] wire113 = wire111 ? wire104 : wire96;
wire [7:0] wire114 = {wire112, wire113};
wire [3:0] wire115 = wire114[7:4];
wire  wire116 = wire97 <= wire103;
wire [3:0] wire117 = wire116 ? wire97 : wire103;
wire [3:0] wire118 = wire116 ? wire103 : wire97;
wire [7:0] wire119 = {wire117, wire118};
wire [3:0] wire120 = wire119[7:4];
wire [7:0] wire121 = {wire112, wire117};
wire [7:0] wire122 = {wire113, wire118};
wire [15:0] wire123 = {wire121, wire122};
wire [7:0] wire124 = wire123[15:8];
wire [3:0] wire125 = wire121[7:4];
wire  wire126 = wire112 <= wire117;
wire [3:0] wire127 = wire126 ? wire112 : wire117;
wire [3:0] wire128 = wire126 ? wire117 : wire112;
wire [7:0] wire129 = {wire127, wire128};
wire [3:0] wire130 = wire129[7:4];
wire  wire131 = wire113 <= wire118;
wire [3:0] wire132 = wire131 ? wire113 : wire118;
wire [3:0] wire133 = wire131 ? wire118 : wire113;
wire [7:0] wire134 = {wire132, wire133};
wire [3:0] wire135 = wire134[7:4];
wire [15:0] wire136 = {wire129, wire134};
wire [7:0] wire137 = wire136[15:8];
wire [7:0] wire138 = {wire133, wire132};
wire [7:0] wire139 = {wire128, wire127};
wire [15:0] wire140 = {wire138, wire139};
wire [31:0] wire141 = {wire92, wire140};
wire [15:0] wire142 = wire141[31:16];
wire [7:0] wire143 = wire92[15:8];
wire [7:0] wire144 = wire140[15:8];
wire [3:0] wire145 = wire138[7:4];
wire [3:0] wire146 = wire139[7:4];
wire  wire147 = wire83 <= wire133;
wire [3:0] wire148 = wire147 ? wire83 : wire133;
wire [3:0] wire149 = wire147 ? wire133 : wire83;
wire [7:0] wire150 = {wire148, wire149};
wire [3:0] wire151 = wire150[7:4];
wire  wire152 = wire84 <= wire132;
wire [3:0] wire153 = wire152 ? wire84 : wire132;
wire [3:0] wire154 = wire152 ? wire132 : wire84;
wire [7:0] wire155 = {wire153, wire154};
wire [3:0] wire156 = wire155[7:4];
wire [7:0] wire157 = {wire148, wire153};
wire [7:0] wire158 = {wire149, wire154};
wire [15:0] wire159 = {wire157, wire158};
wire [7:0] wire160 = wire159[15:8];
wire  wire161 = wire88 <= wire128;
wire [3:0] wire162 = wire161 ? wire88 : wire128;
wire [3:0] wire163 = wire161 ? wire128 : wire88;
wire [7:0] wire164 = {wire162, wire163};
wire [3:0] wire165 = wire164[7:4];
wire  wire166 = wire89 <= wire127;
wire [3:0] wire167 = wire166 ? wire89 : wire127;
wire [3:0] wire168 = wire166 ? wire127 : wire89;
wire [7:0] wire169 = {wire167, wire168};
wire [3:0] wire170 = wire169[7:4];
wire [7:0] wire171 = {wire162, wire167};
wire [7:0] wire172 = {wire163, wire168};
wire [15:0] wire173 = {wire171, wire172};
wire [7:0] wire174 = wire173[15:8];
wire [15:0] wire175 = {wire157, wire171};
wire [15:0] wire176 = {wire158, wire172};
wire [31:0] wire177 = {wire175, wire176};
wire [15:0] wire178 = wire177[31:16];
wire [7:0] wire179 = wire175[15:8];
wire [3:0] wire180 = wire157[7:4];
wire [3:0] wire181 = wire171[7:4];
wire  wire182 = wire148 <= wire162;
wire [3:0] wire183 = wire182 ? wire148 : wire162;
wire [3:0] wire184 = wire182 ? wire162 : wire148;
wire [7:0] wire185 = {wire183, wire184};
wire [3:0] wire186 = wire185[7:4];
wire  wire187 = wire153 <= wire167;
wire [3:0] wire188 = wire187 ? wire153 : wire167;
wire [3:0] wire189 = wire187 ? wire167 : wire153;
wire [7:0] wire190 = {wire188, wire189};
wire [3:0] wire191 = wire190[7:4];
wire [7:0] wire192 = {wire183, wire188};
wire [7:0] wire193 = {wire184, wire189};
wire [15:0] wire194 = {wire192, wire193};
wire [7:0] wire195 = wire194[15:8];
wire [3:0] wire196 = wire192[7:4];
wire  wire197 = wire183 <= wire188;
wire [3:0] wire198 = wire197 ? wire183 : wire188;
wire [3:0] wire199 = wire197 ? wire188 : wire183;
wire [7:0] wire200 = {wire198, wire199};
wire [3:0] wire201 = wire200[7:4];
wire  wire202 = wire184 <= wire189;
wire [3:0] wire203 = wire202 ? wire184 : wire189;
wire [3:0] wire204 = wire202 ? wire189 : wire184;
wire [7:0] wire205 = {wire203, wire204};
wire [3:0] wire206 = wire205[7:4];
wire [15:0] wire207 = {wire200, wire205};
wire  wire208 = wire149 <= wire163;
wire [3:0] wire209 = wire208 ? wire149 : wire163;
wire [3:0] wire210 = wire208 ? wire163 : wire149;
wire [7:0] wire211 = {wire209, wire210};
wire [3:0] wire212 = wire211[7:4];
wire  wire213 = wire154 <= wire168;
wire [3:0] wire214 = wire213 ? wire154 : wire168;
wire [3:0] wire215 = wire213 ? wire168 : wire154;
wire [7:0] wire216 = {wire214, wire215};
wire [3:0] wire217 = wire216[7:4];
wire [7:0] wire218 = {wire209, wire214};
wire [7:0] wire219 = {wire210, wire215};
wire [15:0] wire220 = {wire218, wire219};
wire [7:0] wire221 = wire220[15:8];
wire [3:0] wire222 = wire218[7:4];
wire  wire223 = wire209 <= wire214;
wire [3:0] wire224 = wire223 ? wire209 : wire214;
wire [3:0] wire225 = wire223 ? wire214 : wire209;
wire [7:0] wire226 = {wire224, wire225};
wire [3:0] wire227 = wire226[7:4];
wire  wire228 = wire210 <= wire215;
wire [3:0] wire229 = wire228 ? wire210 : wire215;
wire [3:0] wire230 = wire228 ? wire215 : wire210;
wire [7:0] wire231 = {wire229, wire230};
wire [3:0] wire232 = wire231[7:4];
wire [15:0] wire233 = {wire226, wire231};
wire [31:0] wire234 = {wire207, wire233};
wire [7:0] wire235 = {wire34, wire36};
wire [3:0] wire236 = wire235[7:4];
wire  wire237 = wire34 <= wire36;
wire [3:0] wire238 = wire237 ? wire34 : wire36;
wire [3:0] wire239 = wire237 ? wire36 : wire34;
wire [7:0] wire240 = {wire238, wire239};
wire [3:0] wire241 = wire240[7:4];
wire [7:0] wire242 = {wire37, wire39};
wire [3:0] wire243 = wire242[7:4];
wire  wire244 = wire37 <= wire39;
wire [3:0] wire245 = wire244 ? wire37 : wire39;
wire [3:0] wire246 = wire244 ? wire39 : wire37;
wire [7:0] wire247 = {wire245, wire246};
wire [3:0] wire248 = wire247[7:4];
wire [7:0] wire249 = {wire246, wire245};
wire [15:0] wire250 = {wire240, wire249};
wire [7:0] wire251 = wire250[15:8];
wire [3:0] wire252 = wire249[7:4];
wire  wire253 = wire238 <= wire246;
wire [3:0] wire254 = wire253 ? wire238 : wire246;
wire [3:0] wire255 = wire253 ? wire246 : wire238;
wire [7:0] wire256 = {wire254, wire255};
wire [3:0] wire257 = wire256[7:4];
wire  wire258 = wire239 <= wire245;
wire [3:0] wire259 = wire258 ? wire239 : wire245;
wire [3:0] wire260 = wire258 ? wire245 : wire239;
wire [7:0] wire261 = {wire259, wire260};
wire [3:0] wire262 = wire261[7:4];
wire [7:0] wire263 = {wire254, wire259};
wire [7:0] wire264 = {wire255, wire260};
wire [15:0] wire265 = {wire263, wire264};
wire [7:0] wire266 = wire265[15:8];
wire [3:0] wire267 = wire263[7:4];
wire  wire268 = wire254 <= wire259;
wire [3:0] wire269 = wire268 ? wire254 : wire259;
wire [3:0] wire270 = wire268 ? wire259 : wire254;
wire [7:0] wire271 = {wire269, wire270};
wire [3:0] wire272 = wire271[7:4];
wire  wire273 = wire255 <= wire260;
wire [3:0] wire274 = wire273 ? wire255 : wire260;
wire [3:0] wire275 = wire273 ? wire260 : wire255;
wire [7:0] wire276 = {wire274, wire275};
wire [3:0] wire277 = wire276[7:4];
wire [15:0] wire278 = {wire271, wire276};
wire [7:0] wire279 = {wire43, wire45};
wire [3:0] wire280 = wire279[7:4];
wire  wire281 = wire43 <= wire45;
wire [3:0] wire282 = wire281 ? wire43 : wire45;
wire [3:0] wire283 = wire281 ? wire45 : wire43;
wire [7:0] wire284 = {wire282, wire283};
wire [3:0] wire285 = wire284[7:4];
wire [7:0] wire286 = {wire46, wire48};
wire [3:0] wire287 = wire286[7:4];
wire  wire288 = wire46 <= wire48;
wire [3:0] wire289 = wire288 ? wire46 : wire48;
wire [3:0] wire290 = wire288 ? wire48 : wire46;
wire [7:0] wire291 = {wire289, wire290};
wire [3:0] wire292 = wire291[7:4];
wire [7:0] wire293 = {wire290, wire289};
wire [15:0] wire294 = {wire284, wire293};
wire [7:0] wire295 = wire294[15:8];
wire [3:0] wire296 = wire293[7:4];
wire  wire297 = wire282 <= wire290;
wire [3:0] wire298 = wire297 ? wire282 : wire290;
wire [3:0] wire299 = wire297 ? wire290 : wire282;
wire [7:0] wire300 = {wire298, wire299};
wire [3:0] wire301 = wire300[7:4];
wire  wire302 = wire283 <= wire289;
wire [3:0] wire303 = wire302 ? wire283 : wire289;
wire [3:0] wire304 = wire302 ? wire289 : wire283;
wire [7:0] wire305 = {wire303, wire304};
wire [3:0] wire306 = wire305[7:4];
wire [7:0] wire307 = {wire298, wire303};
wire [7:0] wire308 = {wire299, wire304};
wire [15:0] wire309 = {wire307, wire308};
wire [7:0] wire310 = wire309[15:8];
wire [3:0] wire311 = wire307[7:4];
wire  wire312 = wire298 <= wire303;
wire [3:0] wire313 = wire312 ? wire298 : wire303;
wire [3:0] wire314 = wire312 ? wire303 : wire298;
wire [7:0] wire315 = {wire313, wire314};
wire [3:0] wire316 = wire315[7:4];
wire  wire317 = wire299 <= wire304;
wire [3:0] wire318 = wire317 ? wire299 : wire304;
wire [3:0] wire319 = wire317 ? wire304 : wire299;
wire [7:0] wire320 = {wire318, wire319};
wire [3:0] wire321 = wire320[7:4];
wire [15:0] wire322 = {wire315, wire320};
wire [7:0] wire323 = wire322[15:8];
wire [7:0] wire324 = {wire319, wire318};
wire [7:0] wire325 = {wire314, wire313};
wire [15:0] wire326 = {wire324, wire325};
wire [31:0] wire327 = {wire278, wire326};
wire [15:0] wire328 = wire327[31:16];
wire [7:0] wire329 = wire278[15:8];
wire [7:0] wire330 = wire326[15:8];
wire [3:0] wire331 = wire324[7:4];
wire [3:0] wire332 = wire325[7:4];
wire  wire333 = wire269 <= wire319;
wire [3:0] wire334 = wire333 ? wire269 : wire319;
wire [3:0] wire335 = wire333 ? wire319 : wire269;
wire [7:0] wire336 = {wire334, wire335};
wire [3:0] wire337 = wire336[7:4];
wire  wire338 = wire270 <= wire318;
wire [3:0] wire339 = wire338 ? wire270 : wire318;
wire [3:0] wire340 = wire338 ? wire318 : wire270;
wire [7:0] wire341 = {wire339, wire340};
wire [3:0] wire342 = wire341[7:4];
wire [7:0] wire343 = {wire334, wire339};
wire [7:0] wire344 = {wire335, wire340};
wire [15:0] wire345 = {wire343, wire344};
wire [7:0] wire346 = wire345[15:8];
wire  wire347 = wire274 <= wire314;
wire [3:0] wire348 = wire347 ? wire274 : wire314;
wire [3:0] wire349 = wire347 ? wire314 : wire274;
wire [7:0] wire350 = {wire348, wire349};
wire [3:0] wire351 = wire350[7:4];
wire  wire352 = wire275 <= wire313;
wire [3:0] wire353 = wire352 ? wire275 : wire313;
wire [3:0] wire354 = wire352 ? wire313 : wire275;
wire [7:0] wire355 = {wire353, wire354};
wire [3:0] wire356 = wire355[7:4];
wire [7:0] wire357 = {wire348, wire353};
wire [7:0] wire358 = {wire349, wire354};
wire [15:0] wire359 = {wire357, wire358};
wire [7:0] wire360 = wire359[15:8];
wire [15:0] wire361 = {wire343, wire357};
wire [15:0] wire362 = {wire344, wire358};
wire [31:0] wire363 = {wire361, wire362};
wire [15:0] wire364 = wire363[31:16];
wire [7:0] wire365 = wire361[15:8];
wire [3:0] wire366 = wire343[7:4];
wire [3:0] wire367 = wire357[7:4];
wire  wire368 = wire334 <= wire348;
wire [3:0] wire369 = wire368 ? wire334 : wire348;
wire [3:0] wire370 = wire368 ? wire348 : wire334;
wire [7:0] wire371 = {wire369, wire370};
wire [3:0] wire372 = wire371[7:4];
wire  wire373 = wire339 <= wire353;
wire [3:0] wire374 = wire373 ? wire339 : wire353;
wire [3:0] wire375 = wire373 ? wire353 : wire339;
wire [7:0] wire376 = {wire374, wire375};
wire [3:0] wire377 = wire376[7:4];
wire [7:0] wire378 = {wire369, wire374};
wire [7:0] wire379 = {wire370, wire375};
wire [15:0] wire380 = {wire378, wire379};
wire [7:0] wire381 = wire380[15:8];
wire [3:0] wire382 = wire378[7:4];
wire  wire383 = wire369 <= wire374;
wire [3:0] wire384 = wire383 ? wire369 : wire374;
wire [3:0] wire385 = wire383 ? wire374 : wire369;
wire [7:0] wire386 = {wire384, wire385};
wire [3:0] wire387 = wire386[7:4];
wire  wire388 = wire370 <= wire375;
wire [3:0] wire389 = wire388 ? wire370 : wire375;
wire [3:0] wire390 = wire388 ? wire375 : wire370;
wire [7:0] wire391 = {wire389, wire390};
wire [3:0] wire392 = wire391[7:4];
wire [15:0] wire393 = {wire386, wire391};
wire  wire394 = wire335 <= wire349;
wire [3:0] wire395 = wire394 ? wire335 : wire349;
wire [3:0] wire396 = wire394 ? wire349 : wire335;
wire [7:0] wire397 = {wire395, wire396};
wire [3:0] wire398 = wire397[7:4];
wire  wire399 = wire340 <= wire354;
wire [3:0] wire400 = wire399 ? wire340 : wire354;
wire [3:0] wire401 = wire399 ? wire354 : wire340;
wire [7:0] wire402 = {wire400, wire401};
wire [3:0] wire403 = wire402[7:4];
wire [7:0] wire404 = {wire395, wire400};
wire [7:0] wire405 = {wire396, wire401};
wire [15:0] wire406 = {wire404, wire405};
wire [7:0] wire407 = wire406[15:8];
wire [3:0] wire408 = wire404[7:4];
wire  wire409 = wire395 <= wire400;
wire [3:0] wire410 = wire409 ? wire395 : wire400;
wire [3:0] wire411 = wire409 ? wire400 : wire395;
wire [7:0] wire412 = {wire410, wire411};
wire [3:0] wire413 = wire412[7:4];
wire  wire414 = wire396 <= wire401;
wire [3:0] wire415 = wire414 ? wire396 : wire401;
wire [3:0] wire416 = wire414 ? wire401 : wire396;
wire [7:0] wire417 = {wire415, wire416};
wire [3:0] wire418 = wire417[7:4];
wire [15:0] wire419 = {wire412, wire417};
wire [31:0] wire420 = {wire393, wire419};
wire [15:0] wire421 = wire420[31:16];
wire [7:0] wire422 = wire393[15:8];
wire [7:0] wire423 = wire419[15:8];
wire [7:0] wire424 = {wire416, wire415};
wire [7:0] wire425 = {wire411, wire410};
wire [15:0] wire426 = {wire424, wire425};
wire [7:0] wire427 = {wire390, wire389};
wire [7:0] wire428 = {wire385, wire384};
wire [15:0] wire429 = {wire427, wire428};
wire [31:0] wire430 = {wire426, wire429};
wire [63:0] wire431 = {wire234, wire430};
wire [31:0] wire432 = wire431[63:32];
wire [15:0] wire433 = wire234[31:16];
wire [7:0] wire434 = wire207[15:8];
wire [7:0] wire435 = wire233[15:8];
wire [15:0] wire436 = wire430[31:16];
wire [7:0] wire437 = wire426[15:8];
wire [3:0] wire438 = wire424[7:4];
wire [3:0] wire439 = wire425[7:4];
wire [7:0] wire440 = wire429[15:8];
wire [3:0] wire441 = wire427[7:4];
wire [3:0] wire442 = wire428[7:4];
wire  wire443 = wire198 <= wire416;
wire [3:0] wire444 = wire443 ? wire198 : wire416;
wire [3:0] wire445 = wire443 ? wire416 : wire198;
wire [7:0] wire446 = {wire444, wire445};
wire [3:0] wire447 = wire446[7:4];
wire  wire448 = wire199 <= wire415;
wire [3:0] wire449 = wire448 ? wire199 : wire415;
wire [3:0] wire450 = wire448 ? wire415 : wire199;
wire [7:0] wire451 = {wire449, wire450};
wire [3:0] wire452 = wire451[7:4];
wire [7:0] wire453 = {wire444, wire449};
wire [7:0] wire454 = {wire445, wire450};
wire [15:0] wire455 = {wire453, wire454};
wire [7:0] wire456 = wire455[15:8];
wire  wire457 = wire203 <= wire411;
wire [3:0] wire458 = wire457 ? wire203 : wire411;
wire [3:0] wire459 = wire457 ? wire411 : wire203;
wire [7:0] wire460 = {wire458, wire459};
wire [3:0] wire461 = wire460[7:4];
wire  wire462 = wire204 <= wire410;
wire [3:0] wire463 = wire462 ? wire204 : wire410;
wire [3:0] wire464 = wire462 ? wire410 : wire204;
wire [7:0] wire465 = {wire463, wire464};
wire [3:0] wire466 = wire465[7:4];
wire [7:0] wire467 = {wire458, wire463};
wire [7:0] wire468 = {wire459, wire464};
wire [15:0] wire469 = {wire467, wire468};
wire [7:0] wire470 = wire469[15:8];
wire [15:0] wire471 = {wire453, wire467};
wire [15:0] wire472 = {wire454, wire468};
wire [31:0] wire473 = {wire471, wire472};
wire [15:0] wire474 = wire473[31:16];
wire  wire475 = wire224 <= wire390;
wire [3:0] wire476 = wire475 ? wire224 : wire390;
wire [3:0] wire477 = wire475 ? wire390 : wire224;
wire [7:0] wire478 = {wire476, wire477};
wire [3:0] wire479 = wire478[7:4];
wire  wire480 = wire225 <= wire389;
wire [3:0] wire481 = wire480 ? wire225 : wire389;
wire [3:0] wire482 = wire480 ? wire389 : wire225;
wire [7:0] wire483 = {wire481, wire482};
wire [3:0] wire484 = wire483[7:4];
wire [7:0] wire485 = {wire476, wire481};
wire [7:0] wire486 = {wire477, wire482};
wire [15:0] wire487 = {wire485, wire486};
wire [7:0] wire488 = wire487[15:8];
wire  wire489 = wire229 <= wire385;
wire [3:0] wire490 = wire489 ? wire229 : wire385;
wire [3:0] wire491 = wire489 ? wire385 : wire229;
wire [7:0] wire492 = {wire490, wire491};
wire [3:0] wire493 = wire492[7:4];
wire  wire494 = wire230 <= wire384;
wire [3:0] wire495 = wire494 ? wire230 : wire384;
wire [3:0] wire496 = wire494 ? wire384 : wire230;
wire [7:0] wire497 = {wire495, wire496};
wire [3:0] wire498 = wire497[7:4];
wire [7:0] wire499 = {wire490, wire495};
wire [7:0] wire500 = {wire491, wire496};
wire [15:0] wire501 = {wire499, wire500};
wire [7:0] wire502 = wire501[15:8];
wire [15:0] wire503 = {wire485, wire499};
wire [15:0] wire504 = {wire486, wire500};
wire [31:0] wire505 = {wire503, wire504};
wire [15:0] wire506 = wire505[31:16];
wire [31:0] wire507 = {wire471, wire503};
wire [31:0] wire508 = {wire472, wire504};
wire [63:0] wire509 = {wire507, wire508};
wire [31:0] wire510 = wire509[63:32];
wire [15:0] wire511 = wire507[31:16];
wire [7:0] wire512 = wire471[15:8];
wire [3:0] wire513 = wire453[7:4];
wire [3:0] wire514 = wire467[7:4];
wire [7:0] wire515 = wire503[15:8];
wire [3:0] wire516 = wire485[7:4];
wire [3:0] wire517 = wire499[7:4];
wire  wire518 = wire444 <= wire476;
wire [3:0] wire519 = wire518 ? wire444 : wire476;
wire [3:0] wire520 = wire518 ? wire476 : wire444;
wire [7:0] wire521 = {wire519, wire520};
wire [3:0] wire522 = wire521[7:4];
wire  wire523 = wire449 <= wire481;
wire [3:0] wire524 = wire523 ? wire449 : wire481;
wire [3:0] wire525 = wire523 ? wire481 : wire449;
wire [7:0] wire526 = {wire524, wire525};
wire [3:0] wire527 = wire526[7:4];
wire [7:0] wire528 = {wire519, wire524};
wire [7:0] wire529 = {wire520, wire525};
wire [15:0] wire530 = {wire528, wire529};
wire [7:0] wire531 = wire530[15:8];
wire  wire532 = wire458 <= wire490;
wire [3:0] wire533 = wire532 ? wire458 : wire490;
wire [3:0] wire534 = wire532 ? wire490 : wire458;
wire [7:0] wire535 = {wire533, wire534};
wire [3:0] wire536 = wire535[7:4];
wire  wire537 = wire463 <= wire495;
wire [3:0] wire538 = wire537 ? wire463 : wire495;
wire [3:0] wire539 = wire537 ? wire495 : wire463;
wire [7:0] wire540 = {wire538, wire539};
wire [3:0] wire541 = wire540[7:4];
wire [7:0] wire542 = {wire533, wire538};
wire [7:0] wire543 = {wire534, wire539};
wire [15:0] wire544 = {wire542, wire543};
wire [7:0] wire545 = wire544[15:8];
wire [15:0] wire546 = {wire528, wire542};
wire [15:0] wire547 = {wire529, wire543};
wire [31:0] wire548 = {wire546, wire547};
wire [15:0] wire549 = wire548[31:16];
wire [7:0] wire550 = wire546[15:8];
wire [3:0] wire551 = wire528[7:4];
wire [3:0] wire552 = wire542[7:4];
wire  wire553 = wire519 <= wire533;
wire [3:0] wire554 = wire553 ? wire519 : wire533;
wire [3:0] wire555 = wire553 ? wire533 : wire519;
wire [7:0] wire556 = {wire554, wire555};
wire [3:0] wire557 = wire556[7:4];
wire  wire558 = wire524 <= wire538;
wire [3:0] wire559 = wire558 ? wire524 : wire538;
wire [3:0] wire560 = wire558 ? wire538 : wire524;
wire [7:0] wire561 = {wire559, wire560};
wire [3:0] wire562 = wire561[7:4];
wire [7:0] wire563 = {wire554, wire559};
wire [7:0] wire564 = {wire555, wire560};
wire [15:0] wire565 = {wire563, wire564};
wire [7:0] wire566 = wire565[15:8];
wire [3:0] wire567 = wire563[7:4];
wire  wire568 = wire554 <= wire559;
wire [3:0] wire569 = wire568 ? wire554 : wire559;
wire [3:0] wire570 = wire568 ? wire559 : wire554;
wire [7:0] wire571 = {wire569, wire570};
wire [3:0] wire572 = wire571[7:4];
wire  wire573 = wire555 <= wire560;
wire [3:0] wire574 = wire573 ? wire555 : wire560;
wire [3:0] wire575 = wire573 ? wire560 : wire555;
wire [7:0] wire576 = {wire574, wire575};
wire [3:0] wire577 = wire576[7:4];
wire [15:0] wire578 = {wire571, wire576};
wire  wire579 = wire520 <= wire534;
wire [3:0] wire580 = wire579 ? wire520 : wire534;
wire [3:0] wire581 = wire579 ? wire534 : wire520;
wire [7:0] wire582 = {wire580, wire581};
wire [3:0] wire583 = wire582[7:4];
wire  wire584 = wire525 <= wire539;
wire [3:0] wire585 = wire584 ? wire525 : wire539;
wire [3:0] wire586 = wire584 ? wire539 : wire525;
wire [7:0] wire587 = {wire585, wire586};
wire [3:0] wire588 = wire587[7:4];
wire [7:0] wire589 = {wire580, wire585};
wire [7:0] wire590 = {wire581, wire586};
wire [15:0] wire591 = {wire589, wire590};
wire [7:0] wire592 = wire591[15:8];
wire [3:0] wire593 = wire589[7:4];
wire  wire594 = wire580 <= wire585;
wire [3:0] wire595 = wire594 ? wire580 : wire585;
wire [3:0] wire596 = wire594 ? wire585 : wire580;
wire [7:0] wire597 = {wire595, wire596};
wire [3:0] wire598 = wire597[7:4];
wire  wire599 = wire581 <= wire586;
wire [3:0] wire600 = wire599 ? wire581 : wire586;
wire [3:0] wire601 = wire599 ? wire586 : wire581;
wire [7:0] wire602 = {wire600, wire601};
wire [3:0] wire603 = wire602[7:4];
wire [15:0] wire604 = {wire597, wire602};
wire [31:0] wire605 = {wire578, wire604};
wire  wire606 = wire445 <= wire477;
wire [3:0] wire607 = wire606 ? wire445 : wire477;
wire [3:0] wire608 = wire606 ? wire477 : wire445;
wire [7:0] wire609 = {wire607, wire608};
wire [3:0] wire610 = wire609[7:4];
wire  wire611 = wire450 <= wire482;
wire [3:0] wire612 = wire611 ? wire450 : wire482;
wire [3:0] wire613 = wire611 ? wire482 : wire450;
wire [7:0] wire614 = {wire612, wire613};
wire [3:0] wire615 = wire614[7:4];
wire [7:0] wire616 = {wire607, wire612};
wire [7:0] wire617 = {wire608, wire613};
wire [15:0] wire618 = {wire616, wire617};
wire [7:0] wire619 = wire618[15:8];
wire  wire620 = wire459 <= wire491;
wire [3:0] wire621 = wire620 ? wire459 : wire491;
wire [3:0] wire622 = wire620 ? wire491 : wire459;
wire [7:0] wire623 = {wire621, wire622};
wire [3:0] wire624 = wire623[7:4];
wire  wire625 = wire464 <= wire496;
wire [3:0] wire626 = wire625 ? wire464 : wire496;
wire [3:0] wire627 = wire625 ? wire496 : wire464;
wire [7:0] wire628 = {wire626, wire627};
wire [3:0] wire629 = wire628[7:4];
wire [7:0] wire630 = {wire621, wire626};
wire [7:0] wire631 = {wire622, wire627};
wire [15:0] wire632 = {wire630, wire631};
wire [7:0] wire633 = wire632[15:8];
wire [15:0] wire634 = {wire616, wire630};
wire [15:0] wire635 = {wire617, wire631};
wire [31:0] wire636 = {wire634, wire635};
wire [15:0] wire637 = wire636[31:16];
wire [7:0] wire638 = wire634[15:8];
wire [3:0] wire639 = wire616[7:4];
wire [3:0] wire640 = wire630[7:4];
wire  wire641 = wire607 <= wire621;
wire [3:0] wire642 = wire641 ? wire607 : wire621;
wire [3:0] wire643 = wire641 ? wire621 : wire607;
wire [7:0] wire644 = {wire642, wire643};
wire [3:0] wire645 = wire644[7:4];
wire  wire646 = wire612 <= wire626;
wire [3:0] wire647 = wire646 ? wire612 : wire626;
wire [3:0] wire648 = wire646 ? wire626 : wire612;
wire [7:0] wire649 = {wire647, wire648};
wire [3:0] wire650 = wire649[7:4];
wire [7:0] wire651 = {wire642, wire647};
wire [7:0] wire652 = {wire643, wire648};
wire [15:0] wire653 = {wire651, wire652};
wire [7:0] wire654 = wire653[15:8];
wire [3:0] wire655 = wire651[7:4];
wire  wire656 = wire642 <= wire647;
wire [3:0] wire657 = wire656 ? wire642 : wire647;
wire [3:0] wire658 = wire656 ? wire647 : wire642;
wire [7:0] wire659 = {wire657, wire658};
wire [3:0] wire660 = wire659[7:4];
wire  wire661 = wire643 <= wire648;
wire [3:0] wire662 = wire661 ? wire643 : wire648;
wire [3:0] wire663 = wire661 ? wire648 : wire643;
wire [7:0] wire664 = {wire662, wire663};
wire [3:0] wire665 = wire664[7:4];
wire [15:0] wire666 = {wire659, wire664};
wire  wire667 = wire608 <= wire622;
wire [3:0] wire668 = wire667 ? wire608 : wire622;
wire [3:0] wire669 = wire667 ? wire622 : wire608;
wire [7:0] wire670 = {wire668, wire669};
wire [3:0] wire671 = wire670[7:4];
wire  wire672 = wire613 <= wire627;
wire [3:0] wire673 = wire672 ? wire613 : wire627;
wire [3:0] wire674 = wire672 ? wire627 : wire613;
wire [7:0] wire675 = {wire673, wire674};
wire [3:0] wire676 = wire675[7:4];
wire [7:0] wire677 = {wire668, wire673};
wire [7:0] wire678 = {wire669, wire674};
wire [15:0] wire679 = {wire677, wire678};
wire [7:0] wire680 = wire679[15:8];
wire [3:0] wire681 = wire677[7:4];
wire  wire682 = wire668 <= wire673;
wire [3:0] wire683 = wire682 ? wire668 : wire673;
wire [3:0] wire684 = wire682 ? wire673 : wire668;
wire [7:0] wire685 = {wire683, wire684};
wire [3:0] wire686 = wire685[7:4];
wire  wire687 = wire669 <= wire674;
wire [3:0] wire688 = wire687 ? wire669 : wire674;
wire [3:0] wire689 = wire687 ? wire674 : wire669;
wire [7:0] wire690 = {wire688, wire689};
wire [3:0] wire691 = wire690[7:4];
wire [15:0] wire692 = {wire685, wire690};
wire [31:0] wire693 = {wire666, wire692};
wire [63:0] wire694 = {wire605, wire693};
// effects 
assign guard = wire1;
assign value = wire694;
always@(posedge clk)
begin
	if(rst_n)
		begin
// reset 
		end
	else
		begin
	if(wire1)
		begin
// put  debug code here (display, stop, ...)
		end
		end
end
endmodule